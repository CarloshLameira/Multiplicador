module ACC(Load, Sh, Ad, Clk, Entradas, Saidas);
	
	input Load, Sh, Ad, Clk;
	input [7:0] Entradas;
	output reg [7:0] Saidas;

endmodule
