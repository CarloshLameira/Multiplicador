module Counter(Load, Clk, K);

	input Load, Clk;
	output K;

endmodule

