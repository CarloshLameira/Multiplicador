module Control(Idle, Done, St, Load, Sh, Ad, Clk, k, M);

	input St,Clk,k,M;
	output Idle, Done, Load, Sh, Ad;

endmodule

